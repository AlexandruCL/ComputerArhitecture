library verilog;
use verilog.vl_types.all;
entity rtu2_p1_tb is
end rtu2_p1_tb;
