module mcb(
  input a,
  input b,
  input z,
  input y,
  input ci,
  output w,
  output co
);



endmodule