module bist(
    input clk, rst,
    output [3:0] q
);

