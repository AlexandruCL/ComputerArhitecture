module cl0(
  input x0,
  output a0,
  output b0
);

  assign a0 = x0;
  assign b0 = 1'd1;
endmodule