library verilog;
use verilog.vl_types.all;
entity grade is
end grade;
