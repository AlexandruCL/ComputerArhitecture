library verilog;
use verilog.vl_types.all;
entity ex1c is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        f3              : out    vl_logic
    );
end ex1c;
