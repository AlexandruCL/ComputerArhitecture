library verilog;
use verilog.vl_types.all;
entity ex1c_tb is
end ex1c_tb;
