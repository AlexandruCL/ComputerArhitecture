library verilog;
use verilog.vl_types.all;
entity comb_tb is
end comb_tb;
