library verilog;
use verilog.vl_types.all;
entity prenc_tb is
end prenc_tb;
