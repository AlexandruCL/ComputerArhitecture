library verilog;
use verilog.vl_types.all;
entity c1_add4b_tb is
end c1_add4b_tb;
